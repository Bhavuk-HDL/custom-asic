`default_nettype none

`timescale 10 ns / 1 ps

module codes(
	output wire [31:0]	instruction,
	input wire [7:0]	address
	);

	reg [31:0] instrs [58-1:0];
	
	initial begin
		instrs[0] =  {12'b10101, 5'd0, 3'b000, 5'd1, 7'b0010011}; 
		instrs[1] =  {12'b111, 5'd0, 3'b000, 5'd2, 7'b0010011}; 
		instrs[2] =  {12'b111111111100, 5'd0, 3'b000, 5'd3, 7'b0010011}; 
		instrs[3] =  {12'b1011100, 5'd1, 3'b111, 5'd5, 7'b0010011}; 
		instrs[4] =  {12'b10101, 5'd5, 3'b100, 5'd5, 7'b0010011}; 
		instrs[5] =  {12'b1011100, 5'd1, 3'b110, 5'd6, 7'b0010011}; 
		instrs[6] =  {12'b1011100, 5'd6, 3'b100, 5'd6, 7'b0010011}; 
		instrs[7] =  {12'b111, 5'd1, 3'b000, 5'd7, 7'b0010011}; 
		instrs[8] =  {12'b11101, 5'd7, 3'b100, 5'd7, 7'b0010011}; 
		instrs[9] =  {6'b000000, 6'b110, 5'd1, 3'b001, 5'd8, 7'b0010011}; 
		instrs[10] = {12'b10101000001, 5'd8, 3'b100, 5'd8, 7'b0010011}; 
		instrs[11] = {6'b000000, 6'b10, 5'd1, 3'b101, 5'd9, 7'b0010011}; 
		instrs[12] = {12'b100, 5'd9, 3'b100, 5'd9, 7'b0010011}; 
		instrs[13] = {7'b0000000, 5'd2, 5'd1, 3'b111, 5'd10, 7'b0110011}; 
		instrs[14] = {12'b100, 5'd10, 3'b100, 5'd10, 7'b0010011}; 
		instrs[15] = {7'b0000000, 5'd2, 5'd1, 3'b110, 5'd11, 7'b0110011}; 
		instrs[16] = {12'b10110, 5'd11, 3'b100, 5'd11, 7'b0010011}; 
		instrs[17] = {7'b0000000, 5'd2, 5'd1, 3'b100, 5'd12, 7'b0110011}; 
		instrs[18] = {12'b10011, 5'd12, 3'b100, 5'd12, 7'b0010011}; 
		instrs[19] = {7'b0000000, 5'd2, 5'd1, 3'b000, 5'd13, 7'b0110011}; 
		instrs[20] = {12'b11101, 5'd13, 3'b100, 5'd13, 7'b0010011}; 
		instrs[21] = {7'b0100000, 5'd2, 5'd1, 3'b000, 5'd14, 7'b0110011}; 
		instrs[22] = {12'b1111, 5'd14, 3'b100, 5'd14, 7'b0010011}; 
		instrs[23] = {7'b0000000, 5'd2, 5'd2, 3'b001, 5'd15, 7'b0110011}; 
		instrs[24] = {12'b1110000001, 5'd15, 3'b100, 5'd15, 7'b0010011}; 
		instrs[25] = {7'b0000000, 5'd2, 5'd1, 3'b101, 5'd16, 7'b0110011}; 
		instrs[26] = {12'b1, 5'd16, 3'b100, 5'd16, 7'b0010011}; 
		instrs[27] = {7'b0000000, 5'd1, 5'd2, 3'b011, 5'd17, 7'b0110011}; 
		instrs[28] = {12'b0, 5'd17, 3'b100, 5'd17, 7'b0010011}; 
		instrs[29] = {12'b10101, 5'd2, 3'b011, 5'd18, 7'b0010011}; 
		instrs[30] = {12'b0, 5'd18, 3'b100, 5'd18, 7'b0010011}; 
		instrs[31] = {20'b00000000000000000000, 5'd19, 7'b0110111}; 
		instrs[32] = {12'b1, 5'd19, 3'b100, 5'd19, 7'b0010011}; 
		instrs[33] = {6'b010000, 6'b1, 5'd3, 3'b101, 5'd20, 7'b0010011}; 
		instrs[34] = {12'b111111111111, 5'd20, 3'b100, 5'd20, 7'b0010011}; 
		instrs[35] = {7'b0000000, 5'd1, 5'd3, 3'b010, 5'd21, 7'b0110011}; 
		instrs[36] = {12'b0, 5'd21, 3'b100, 5'd21, 7'b0010011}; 
		instrs[37] = {12'b1, 5'd3, 3'b010, 5'd22, 7'b0010011}; 
		instrs[38] = {12'b0, 5'd22, 3'b100, 5'd22, 7'b0010011}; 
		instrs[39] = {7'b0100000, 5'd2, 5'd1, 3'b101, 5'd23, 7'b0110011}; 
		instrs[40] = {12'b1, 5'd23, 3'b100, 5'd23, 7'b0010011}; 
		instrs[41] = {20'b00000000000000000100, 5'd4, 7'b0010111}; 
		instrs[42] = {6'b000000, 6'b111, 5'd4, 3'b101, 5'd24, 7'b0010011}; 
		instrs[43] = {12'b10000000, 5'd24, 3'b100, 5'd24, 7'b0010011}; 
		instrs[44] = {1'b0, 10'b0000000010, 1'b0, 8'b00000000, 5'd25, 7'b1101111}; 
		instrs[45] = {20'b00000000000000000000, 5'd4, 7'b0010111}; 
		instrs[46] = {7'b0000000, 5'd4, 5'd25, 3'b100, 5'd25, 7'b0110011}; 
		instrs[47] = {12'b1, 5'd25, 3'b100, 5'd25, 7'b0010011}; 
		instrs[48] = {12'b10000, 5'd4, 3'b000, 5'd26, 7'b1100111}; 
		instrs[49] = {7'b0100000, 5'd4, 5'd26, 3'b000, 5'd26, 7'b0110011}; 
		instrs[50] = {12'b111111110001, 5'd26, 3'b000, 5'd26, 7'b0010011}; 
		instrs[51] = {7'b0000000, 5'd1, 5'd2, 3'b010, 5'b00001, 7'b0100011}; 
		instrs[52] = {12'b1, 5'd2, 3'b010, 5'd27, 7'b0000011}; 
		instrs[53] = {12'b10100, 5'd27, 3'b100, 5'd27, 7'b0010011}; 
		instrs[54] = {12'b1, 5'd0, 3'b000, 5'd28, 7'b0010011}; 
		instrs[55] = {12'b1, 5'd0, 3'b000, 5'd29, 7'b0010011}; 
		instrs[56] = {12'b1, 5'd0, 3'b000, 5'd30, 7'b0010011}; 
		instrs[57] = {1'b0, 10'b0000000000, 1'b0, 8'b00000000, 5'd0, 7'b1101111};
	end
	
	assign instruction = instrs[address];
	
endmodule

`default_nettype wire
